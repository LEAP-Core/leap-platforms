interface ChannelIO;
endinterface

module mkChannelIO(ChannelIO);
endmodule
