
interface TopLevelWires;
endinterface

interface TopLevelWiresDriver;

    interface TopLevelWires wires_out;

endinterface

module mkTopLevelWiresDriver (TopLevelWiresDriver);

    interface TopLevelWires wires_out;
    endinterface

endmodule
