import channelio::*;

interface RRRClient;
endinterface

module mkRRRClient#(ChannelIO channel) (RRRClient);
endmodule
