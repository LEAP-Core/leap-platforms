// Simulation Physical Platform

`include "unix_pipe_device.bsh"

// PHYSICAL_DRIVERS

// This represents the collection of all platform capabilities which the
// rest of the FPGA uses to interact with the outside world.
// We use other modules to actually do the work.

interface PHYSICAL_DRIVERS;

    interface UNIX_PIPE_DRIVER unixPipeDriver;

    // each set of physical drivers must support a soft reset method
    method Action soft_reset();

endinterface

// TOP_LEVEL_WIRES

// The TOP_LEVEL_WIRES is the datatype which gets passed to the top level
// and output as input/output wires. These wires are then connected to
// physical pins on the FPGA as specified in the accompanying UCF file.
// These wires are defined in the individual devices.

interface TOP_LEVEL_WIRES;

    interface UNIX_PIPE_WIRES unixPipeWires;
    
endinterface

// PHYSICAL_PLATFORM

// The platform is the aggregation of wires and drivers.

interface PHYSICAL_PLATFORM;

    interface PHYSICAL_DRIVERS physicalDrivers;
    interface TOP_LEVEL_WIRES  topLevelWires;

endinterface

// mkPhysicalPlatform

// This is a convenient way for the outside world to instantiate all the devices
// and an aggregation of all the wires.

module mkPhysicalPlatform
       //interface: 
                    (PHYSICAL_PLATFORM);
    
    // Submodules
    
    UNIX_PIPE_DEVICE unix_pipe_device  <- mkUNIXPipeDevice();
    
    // Aggregate the drivers
    
    interface PHYSICAL_DRIVERS physicalDrivers;
    
        interface unixPipeDriver = unix_pipe_device.driver;

        // Soft Reset
        method Action soft_reset() if (unix_pipe_device.driver.soft_reset_requested());
            unix_pipe_device.driver.soft_reset_received();
        endmethod

    endinterface
    
    // Aggregate the wires
    
    interface TOP_LEVEL_WIRES topLevelWires;
    
        interface unixPipeWires  = unix_pipe_device.wires;

    endinterface
               
endmodule
