`include "physical_platform.bsh"

interface CHANNEL_IO;
endinterface

module mkChannelIO#(PHYSICAL_DRIVERS drivers) (CHANNEL_IO);
endmodule
