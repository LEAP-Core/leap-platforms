//
// Copyright (C) 2008 Intel Corporation
//
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
//

//
// Instantiate Clock Buffers for DCM/PLL inputs and outputs
//

import Clocks::*;

//
// General interface that wraps a clock
//

interface CLOCK_WRAPPER_IFC;
    
    interface Clock clock;
    
endinterface

//
// Clock Buffer
//

// import the verilog
import "BVI"
module clock_buffer#(Clock inputClock)
    // interface:
        (CLOCK_WRAPPER_IFC);

    input_clock (CLK_IN) = inputClock;
    
    output_clock clock (CLK_OUT);

endmodule

// wrap it in a nicer module
module mkClockBuffer#(Clock inputClock)
    // interface:
        (Clock);
    
    let buffer <- clock_buffer(inputClock);
    
    return buffer.clock;
    
endmodule

//
// Clock Input Buffer
//

// import the verilog
import "BVI"
module clock_input_buffer#(Clock inputClock)
    // interface:
        (CLOCK_WRAPPER_IFC);

    input_clock (CLK_IN) = inputClock;
    
    output_clock clock (CLK_OUT);

endmodule

// wrap it in a nicer module
module mkClockInputBuffer#(Clock inputClock)
    // interface:
        (Clock);
    
    let buffer <- clock_input_buffer(inputClock);
    
    return buffer.clock;
    
endmodule
