import low_level_platform_interface::*;

interface Memory;
endinterface

module mkMemory#(LowLevelPlatformInterface llpint) (Memory);
endmodule
