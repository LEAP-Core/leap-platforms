import rrr::*;
import toplevel_wires::*;

interface Memory;
endinterface

module mkMemory#(RPCClient rpcClient, TopLevelWiresDriver wires) (Memory);
endmodule
