`include "toplevel_wires.bsh"

interface ChannelIO;
endinterface

module mkChannelIO#(TopLevelWiresDriver wires) (ChannelIO);
endmodule
