`include "physical_platform.bsh"

interface ChannelIO;
endinterface

module mkChannelIO#(PHYSICAL_DRIVERS drivers) (ChannelIO);
endmodule
