//
// Copyright (c) 2015, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//


//
// mkLEAPCrossingReg --
//   A wrapper for Bluespec's mkNullCrossingReg, which allows us to make 
//   timing assertions during physical synthesis.  
// 

import "BVI" leap_crossing_reg = module mkLEAPCrossingReg#(Clock dstClock, t_REG initialValue)
    // interface:
    (CrossingReg#(t_REG))

    // provisos
    provisos(Bits#(t_REG, t_REG_SZ));

    parameter INITIAL_VALUE = pack(initialValue);
    parameter WIDTH = valueof(t_REG_SZ);

    default_reset rst (RST_N);
    default_clock clk (CLK);
    
    input_clock dstClockIn (CLK_DST)  = dstClock;

    method readData _read();
    method readDataCrossed crossed() clocked_by(dstClockIn);
    method _write(writeData) enable(writeEnable);

    schedule _write C _write;
    schedule (crossed, _read) CF (crossed, _read);
    schedule (_read) SB _write;

endmodule