`include "asim/provides/low_level_platform_interface.bsh"


interface VIRTUAL_DEVICES;

endinterface

module mkVirtualDevices#(LowLevelPlatformInterface llpint) (VIRTUAL_DEVICES);

endmodule
