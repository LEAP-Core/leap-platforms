//
// Copyright (C) 2009 Intel Corporation
//
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
//

//
// Common definition of the interface to a scratchpad virtual device.
//

//
// Interface to a single scratchpad port.  By having separate ports defined
// for each scratchpad, instead of adding a port argument to the methods,
// this module is capable of defining the relative priority of the ports.
//
interface SCRATCHPAD_MEMORY_PORT;
    interface MEMORY_IFC#(SCRATCHPAD_MEM_ADDRESS, SCRATCHPAD_MEM_VALUE) mem;

    // Initialize a port, requesting an allocation of allocLastWordIdx + 1
    // SCRATCHPAD_MEM_VALUE sized words.
    method ActionValue#(Bool) init(SCRATCHPAD_MEM_ADDRESS allocLastWordIdx);
endinterface: SCRATCHPAD_MEMORY_PORT

//
// A scratchpad interface has one memory interface for each client.  Using
// a vector of MEMORY_IFCs instead of adding a port parameter to a
// MEMORY_IFC-like interface makes the scratchpad interchangeable with
// other memories in the clients.
//
interface SCRATCHPAD_MEMORY_VIRTUAL_DEVICE;
    interface Vector#(SCRATCHPAD_N_CLIENTS, SCRATCHPAD_MEMORY_PORT) ports;
endinterface: SCRATCHPAD_MEMORY_VIRTUAL_DEVICE
