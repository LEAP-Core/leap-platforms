import channelio::*;

interface RPCClient;
endinterface

module mkRPCClient#(ChannelIO channel) (RPCClient);
endmodule
