
module clock_import(clk_in,
		    clk_out);
   input clk_in;
   output clk_out;

   assign clk_out = clk_in;
   
endmodule